`timescale 1ns / 1ps

module imm_Gen (
    input  logic [31:0] inst_code,
    output logic [31:0] Imm_out
);

  // falta implementar o I_TYPE do inst_code para o Opcode 0010011
  always_comb
    case (inst_code[6:0])
      7'b0010011: //I_TYPE
      Imm_out = {inst_code[31] ? 20'hFFFFF : 20'b0, inst_code[31:20]};

      7'b0000011:  /*I-type load part*/
      Imm_out = {inst_code[31] ? 20'hFFFFF : 20'b0, inst_code[31:20]};

      7'b0100011:  /*S-type*/
      Imm_out = {inst_code[31] ? 20'hFFFFF : 20'b0, inst_code[31:25], inst_code[11:7]};

      7'b1100011:  /*B-type*/
      Imm_out = {
        inst_code[31] ? 19'h7FFFF : 19'b0,
        inst_code[31],
        inst_code[7],
        inst_code[30:25],
        inst_code[11:8],
        1'b0
      };

      7'b1101111:  /*J-type*/
      Imm_out = {
        inst_code[31] ? 11'b1 : 11'b0, // 20 bits
        inst_code[31:12],
        1'b0
      };
      //$signed(

      7'b1100111:  /*I-type jalr part*/
      Imm_out = {inst_code[31] ? 20'hFFFFF : 20'b0, inst_code[31:20]};

      default: Imm_out = {32'b0};

    endcase
    // JAL : JAL rd, i -> 20bits portanto, rd = PC + 4 e PC = PC + i;
    // JALR: JALR xn, xm, i -> 12bits portanto, xn = PC + 4 e  PC = xm + i;

endmodule
